-- PongFPGA.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PongFPGA is
	port (
		clk_clk          : in  std_logic                    := '0'; --   clk.clk
		hdmi_output_clk  : out std_logic;                           --  hdmi.output_clk
		hdmi_output_data : out std_logic_vector(2 downto 0);        --      .output_data
		reset_reset_n    : in  std_logic                    := '0'  -- reset.reset_n
	);
end entity PongFPGA;

architecture rtl of PongFPGA is
	component AvalonRAMConnector is
		generic (
			DISPLAY_RES_WIDTH  : integer := 640;
			DISPLAY_RES_HEIGHT : integer := 480;
			PX_X_SPLIT         : integer := 20;
			PX_Y_SPLIT         : integer := 20
		);
		port (
			address   : out std_logic_vector(20 downto 0);                    -- address
			read      : out std_logic;                                        -- read
			readdata  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			write     : out std_logic;                                        -- write
			writedata : out std_logic_vector(7 downto 0);                     -- writedata
			px_clk    : in  std_logic                     := 'X';             -- clk
			px_x      : in  std_logic_vector(11 downto 0) := (others => 'X'); -- px_x
			px_y      : in  std_logic_vector(11 downto 0) := (others => 'X'); -- px_y
			px_color  : out std_logic;                                        -- px_color
			reset     : in  std_logic                     := 'X'              -- reset
		);
	end component AvalonRAMConnector;

	component HDMIDriver is
		generic (
			DISPLAY_RES_WIDTH  : integer := 640;
			DISPLAY_RES_HEIGHT : integer := 480;
			PX_FRONT_PORCH     : integer := 16;
			PX_SYNC_PULSE      : integer := 96;
			PX_BACK_PORCH      : integer := 48;
			ROW_FRONT_PORCH    : integer := 10;
			ROW_SYNC_PULSE     : integer := 2;
			ROW_BACK_PORCH     : integer := 33
		);
		port (
			px_clk      : in  std_logic                     := 'X'; -- clk
			px_x        : out std_logic_vector(11 downto 0);        -- px_x
			px_y        : out std_logic_vector(11 downto 0);        -- px_y
			px_color    : in  std_logic                     := 'X'; -- px_color
			bit_clk     : in  std_logic                     := 'X'; -- clk
			output_clk  : out std_logic;                            -- output_clk
			output_data : out std_logic_vector(2 downto 0)          -- output_data
		);
	end component HDMIDriver;

	component PongFPGA_NIOS is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(12 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(11 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component PongFPGA_NIOS;

	component PongFPGA_PLL is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component PongFPGA_PLL;

	component PongFPGA_VRAM is
		port (
			clk         : in  std_logic                    := 'X';             -- clk
			address     : in  std_logic_vector(6 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                    := 'X';             -- clken
			chipselect  : in  std_logic                    := 'X';             -- chipselect
			write       : in  std_logic                    := 'X';             -- write
			readdata    : out std_logic_vector(7 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			reset       : in  std_logic                    := 'X';             -- reset
			reset_req   : in  std_logic                    := 'X';             -- reset_req
			address2    : in  std_logic_vector(6 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                    := 'X';             -- chipselect
			clken2      : in  std_logic                    := 'X';             -- clken
			write2      : in  std_logic                    := 'X';             -- write
			readdata2   : out std_logic_vector(7 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			clk2        : in  std_logic                    := 'X';             -- clk
			reset2      : in  std_logic                    := 'X';             -- reset
			reset_req2  : in  std_logic                    := 'X';             -- reset_req
			freeze      : in  std_logic                    := 'X'              -- freeze
		);
	end component PongFPGA_VRAM;

	component PongFPGA_mm_interconnect_0 is
		port (
			PLL_c1_clk                                                     : in  std_logic                     := 'X';             -- clk
			AvalonRAMConnector_mono_1b_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			AvalonRAMConnector_mono_1b_0_avalon_master_address             : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			AvalonRAMConnector_mono_1b_0_avalon_master_read                : in  std_logic                     := 'X';             -- read
			AvalonRAMConnector_mono_1b_0_avalon_master_readdata            : out std_logic_vector(7 downto 0);                     -- readdata
			AvalonRAMConnector_mono_1b_0_avalon_master_write               : in  std_logic                     := 'X';             -- write
			AvalonRAMConnector_mono_1b_0_avalon_master_writedata           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			VRAM_s2_address                                                : out std_logic_vector(6 downto 0);                     -- address
			VRAM_s2_write                                                  : out std_logic;                                        -- write
			VRAM_s2_readdata                                               : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			VRAM_s2_writedata                                              : out std_logic_vector(7 downto 0);                     -- writedata
			VRAM_s2_chipselect                                             : out std_logic;                                        -- chipselect
			VRAM_s2_clken                                                  : out std_logic                                         -- clken
		);
	end component PongFPGA_mm_interconnect_0;

	component PongFPGA_mm_interconnect_1 is
		port (
			CLK_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			PLL_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			NIOS_reset_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			PLL_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			NIOS_data_master_address                              : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			NIOS_data_master_waitrequest                          : out std_logic;                                        -- waitrequest
			NIOS_data_master_byteenable                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS_data_master_read                                 : in  std_logic                     := 'X';             -- read
			NIOS_data_master_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS_data_master_write                                : in  std_logic                     := 'X';             -- write
			NIOS_data_master_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS_data_master_debugaccess                          : in  std_logic                     := 'X';             -- debugaccess
			NIOS_instruction_master_address                       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			NIOS_instruction_master_waitrequest                   : out std_logic;                                        -- waitrequest
			NIOS_instruction_master_read                          : in  std_logic                     := 'X';             -- read
			NIOS_instruction_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS_debug_mem_slave_address                          : out std_logic_vector(8 downto 0);                     -- address
			NIOS_debug_mem_slave_write                            : out std_logic;                                        -- write
			NIOS_debug_mem_slave_read                             : out std_logic;                                        -- read
			NIOS_debug_mem_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS_debug_mem_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS_debug_mem_slave_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS_debug_mem_slave_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			NIOS_debug_mem_slave_debugaccess                      : out std_logic;                                        -- debugaccess
			PLL_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			PLL_pll_slave_write                                   : out std_logic;                                        -- write
			PLL_pll_slave_read                                    : out std_logic;                                        -- read
			PLL_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLL_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			VRAM_s1_address                                       : out std_logic_vector(6 downto 0);                     -- address
			VRAM_s1_write                                         : out std_logic;                                        -- write
			VRAM_s1_readdata                                      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			VRAM_s1_writedata                                     : out std_logic_vector(7 downto 0);                     -- writedata
			VRAM_s1_chipselect                                    : out std_logic;                                        -- chipselect
			VRAM_s1_clken                                         : out std_logic                                         -- clken
		);
	end component PongFPGA_mm_interconnect_1;

	component PongFPGA_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component PongFPGA_irq_mapper;

	component pongfpga_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component pongfpga_rst_controller;

	component pongfpga_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component pongfpga_rst_controller_002;

	signal pll_c0_clk                                           : std_logic;                     -- PLL:c0 -> [NIOS:clk, VRAM:clk, irq_mapper:clk, mm_interconnect_1:PLL_c0_clk, rst_controller_001:clk]
	signal pll_c1_clk                                           : std_logic;                     -- PLL:c1 -> [AvalonRAMConnector_mono_1b_0:px_clk, HDMIDriver_mono_1b_0:px_clk, VRAM:clk2, mm_interconnect_0:PLL_c1_clk, rst_controller:clk]
	signal pll_c2_clk                                           : std_logic;                     -- PLL:c2 -> HDMIDriver_mono_1b_0:bit_clk
	signal hdmidriver_mono_1b_0_px_address_px_x                 : std_logic_vector(11 downto 0); -- HDMIDriver_mono_1b_0:px_x -> AvalonRAMConnector_mono_1b_0:px_x
	signal hdmidriver_mono_1b_0_px_address_px_y                 : std_logic_vector(11 downto 0); -- HDMIDriver_mono_1b_0:px_y -> AvalonRAMConnector_mono_1b_0:px_y
	signal avalonramconnector_mono_1b_0_px_color_px_color       : std_logic;                     -- AvalonRAMConnector_mono_1b_0:px_color -> HDMIDriver_mono_1b_0:px_color
	signal avalonramconnector_mono_1b_0_avalon_master_readdata  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:AvalonRAMConnector_mono_1b_0_avalon_master_readdata -> AvalonRAMConnector_mono_1b_0:readdata
	signal avalonramconnector_mono_1b_0_avalon_master_address   : std_logic_vector(20 downto 0); -- AvalonRAMConnector_mono_1b_0:address -> mm_interconnect_0:AvalonRAMConnector_mono_1b_0_avalon_master_address
	signal avalonramconnector_mono_1b_0_avalon_master_read      : std_logic;                     -- AvalonRAMConnector_mono_1b_0:read -> mm_interconnect_0:AvalonRAMConnector_mono_1b_0_avalon_master_read
	signal avalonramconnector_mono_1b_0_avalon_master_write     : std_logic;                     -- AvalonRAMConnector_mono_1b_0:write -> mm_interconnect_0:AvalonRAMConnector_mono_1b_0_avalon_master_write
	signal avalonramconnector_mono_1b_0_avalon_master_writedata : std_logic_vector(7 downto 0);  -- AvalonRAMConnector_mono_1b_0:writedata -> mm_interconnect_0:AvalonRAMConnector_mono_1b_0_avalon_master_writedata
	signal mm_interconnect_0_vram_s2_chipselect                 : std_logic;                     -- mm_interconnect_0:VRAM_s2_chipselect -> VRAM:chipselect2
	signal mm_interconnect_0_vram_s2_readdata                   : std_logic_vector(7 downto 0);  -- VRAM:readdata2 -> mm_interconnect_0:VRAM_s2_readdata
	signal mm_interconnect_0_vram_s2_address                    : std_logic_vector(6 downto 0);  -- mm_interconnect_0:VRAM_s2_address -> VRAM:address2
	signal mm_interconnect_0_vram_s2_write                      : std_logic;                     -- mm_interconnect_0:VRAM_s2_write -> VRAM:write2
	signal mm_interconnect_0_vram_s2_writedata                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:VRAM_s2_writedata -> VRAM:writedata2
	signal mm_interconnect_0_vram_s2_clken                      : std_logic;                     -- mm_interconnect_0:VRAM_s2_clken -> VRAM:clken2
	signal nios_data_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_1:NIOS_data_master_readdata -> NIOS:d_readdata
	signal nios_data_master_waitrequest                         : std_logic;                     -- mm_interconnect_1:NIOS_data_master_waitrequest -> NIOS:d_waitrequest
	signal nios_data_master_debugaccess                         : std_logic;                     -- NIOS:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:NIOS_data_master_debugaccess
	signal nios_data_master_address                             : std_logic_vector(12 downto 0); -- NIOS:d_address -> mm_interconnect_1:NIOS_data_master_address
	signal nios_data_master_byteenable                          : std_logic_vector(3 downto 0);  -- NIOS:d_byteenable -> mm_interconnect_1:NIOS_data_master_byteenable
	signal nios_data_master_read                                : std_logic;                     -- NIOS:d_read -> mm_interconnect_1:NIOS_data_master_read
	signal nios_data_master_write                               : std_logic;                     -- NIOS:d_write -> mm_interconnect_1:NIOS_data_master_write
	signal nios_data_master_writedata                           : std_logic_vector(31 downto 0); -- NIOS:d_writedata -> mm_interconnect_1:NIOS_data_master_writedata
	signal nios_instruction_master_readdata                     : std_logic_vector(31 downto 0); -- mm_interconnect_1:NIOS_instruction_master_readdata -> NIOS:i_readdata
	signal nios_instruction_master_waitrequest                  : std_logic;                     -- mm_interconnect_1:NIOS_instruction_master_waitrequest -> NIOS:i_waitrequest
	signal nios_instruction_master_address                      : std_logic_vector(11 downto 0); -- NIOS:i_address -> mm_interconnect_1:NIOS_instruction_master_address
	signal nios_instruction_master_read                         : std_logic;                     -- NIOS:i_read -> mm_interconnect_1:NIOS_instruction_master_read
	signal mm_interconnect_1_nios_debug_mem_slave_readdata      : std_logic_vector(31 downto 0); -- NIOS:debug_mem_slave_readdata -> mm_interconnect_1:NIOS_debug_mem_slave_readdata
	signal mm_interconnect_1_nios_debug_mem_slave_waitrequest   : std_logic;                     -- NIOS:debug_mem_slave_waitrequest -> mm_interconnect_1:NIOS_debug_mem_slave_waitrequest
	signal mm_interconnect_1_nios_debug_mem_slave_debugaccess   : std_logic;                     -- mm_interconnect_1:NIOS_debug_mem_slave_debugaccess -> NIOS:debug_mem_slave_debugaccess
	signal mm_interconnect_1_nios_debug_mem_slave_address       : std_logic_vector(8 downto 0);  -- mm_interconnect_1:NIOS_debug_mem_slave_address -> NIOS:debug_mem_slave_address
	signal mm_interconnect_1_nios_debug_mem_slave_read          : std_logic;                     -- mm_interconnect_1:NIOS_debug_mem_slave_read -> NIOS:debug_mem_slave_read
	signal mm_interconnect_1_nios_debug_mem_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_1:NIOS_debug_mem_slave_byteenable -> NIOS:debug_mem_slave_byteenable
	signal mm_interconnect_1_nios_debug_mem_slave_write         : std_logic;                     -- mm_interconnect_1:NIOS_debug_mem_slave_write -> NIOS:debug_mem_slave_write
	signal mm_interconnect_1_nios_debug_mem_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_1:NIOS_debug_mem_slave_writedata -> NIOS:debug_mem_slave_writedata
	signal mm_interconnect_1_pll_pll_slave_readdata             : std_logic_vector(31 downto 0); -- PLL:readdata -> mm_interconnect_1:PLL_pll_slave_readdata
	signal mm_interconnect_1_pll_pll_slave_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_1:PLL_pll_slave_address -> PLL:address
	signal mm_interconnect_1_pll_pll_slave_read                 : std_logic;                     -- mm_interconnect_1:PLL_pll_slave_read -> PLL:read
	signal mm_interconnect_1_pll_pll_slave_write                : std_logic;                     -- mm_interconnect_1:PLL_pll_slave_write -> PLL:write
	signal mm_interconnect_1_pll_pll_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_1:PLL_pll_slave_writedata -> PLL:writedata
	signal mm_interconnect_1_vram_s1_chipselect                 : std_logic;                     -- mm_interconnect_1:VRAM_s1_chipselect -> VRAM:chipselect
	signal mm_interconnect_1_vram_s1_readdata                   : std_logic_vector(7 downto 0);  -- VRAM:readdata -> mm_interconnect_1:VRAM_s1_readdata
	signal mm_interconnect_1_vram_s1_address                    : std_logic_vector(6 downto 0);  -- mm_interconnect_1:VRAM_s1_address -> VRAM:address
	signal mm_interconnect_1_vram_s1_write                      : std_logic;                     -- mm_interconnect_1:VRAM_s1_write -> VRAM:write
	signal mm_interconnect_1_vram_s1_writedata                  : std_logic_vector(7 downto 0);  -- mm_interconnect_1:VRAM_s1_writedata -> VRAM:writedata
	signal mm_interconnect_1_vram_s1_clken                      : std_logic;                     -- mm_interconnect_1:VRAM_s1_clken -> VRAM:clken
	signal nios_irq_irq                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOS:irq
	signal rst_controller_reset_out_reset                       : std_logic;                     -- rst_controller:reset_out -> [AvalonRAMConnector_mono_1b_0:reset, VRAM:reset2, mm_interconnect_0:AvalonRAMConnector_mono_1b_0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_reset_out_reset_req                   : std_logic;                     -- rst_controller:reset_req -> [VRAM:reset_req2, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                   : std_logic;                     -- rst_controller_001:reset_out -> [VRAM:reset, irq_mapper:reset, mm_interconnect_1:NIOS_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req               : std_logic;                     -- rst_controller_001:reset_req -> [NIOS:reset_req, VRAM:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_002_reset_out_reset                   : std_logic;                     -- rst_controller_002:reset_out -> [PLL:reset, mm_interconnect_1:PLL_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                              : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv         : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> NIOS:reset_n

begin

	avalonramconnector_mono_1b_0 : component AvalonRAMConnector
		generic map (
			DISPLAY_RES_WIDTH  => 640,
			DISPLAY_RES_HEIGHT => 480,
			PX_X_SPLIT         => 20,
			PX_Y_SPLIT         => 20
		)
		port map (
			address   => avalonramconnector_mono_1b_0_avalon_master_address,   -- avalon_master.address
			read      => avalonramconnector_mono_1b_0_avalon_master_read,      --              .read
			readdata  => avalonramconnector_mono_1b_0_avalon_master_readdata,  --              .readdata
			write     => avalonramconnector_mono_1b_0_avalon_master_write,     --              .write
			writedata => avalonramconnector_mono_1b_0_avalon_master_writedata, --              .writedata
			px_clk    => pll_c1_clk,                                           --        px_clk.clk
			px_x      => hdmidriver_mono_1b_0_px_address_px_x,                 --    px_address.px_x
			px_y      => hdmidriver_mono_1b_0_px_address_px_y,                 --              .px_y
			px_color  => avalonramconnector_mono_1b_0_px_color_px_color,       --      px_color.px_color
			reset     => rst_controller_reset_out_reset                        --         reset.reset
		);

	hdmidriver_mono_1b_0 : component HDMIDriver
		generic map (
			DISPLAY_RES_WIDTH  => 640,
			DISPLAY_RES_HEIGHT => 480,
			PX_FRONT_PORCH     => 16,
			PX_SYNC_PULSE      => 96,
			PX_BACK_PORCH      => 48,
			ROW_FRONT_PORCH    => 10,
			ROW_SYNC_PULSE     => 2,
			ROW_BACK_PORCH     => 33
		)
		port map (
			px_clk      => pll_c1_clk,                                     --      clock.clk
			px_x        => hdmidriver_mono_1b_0_px_address_px_x,           -- px_address.px_x
			px_y        => hdmidriver_mono_1b_0_px_address_px_y,           --           .px_y
			px_color    => avalonramconnector_mono_1b_0_px_color_px_color, --   px_color.px_color
			bit_clk     => pll_c2_clk,                                     --    bit_clk.clk
			output_clk  => hdmi_output_clk,                                --       hdmi.output_clk
			output_data => hdmi_output_data                                --           .output_data
		);

	nios : component PongFPGA_NIOS
		port map (
			clk                                 => pll_c0_clk,                                         --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,       --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,             --                          .reset_req
			d_address                           => nios_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_data_master_read,                              --                          .read
			d_readdata                          => nios_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_data_master_write,                             --                          .write
			d_writedata                         => nios_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_instruction_master_read,                       --                          .read
			i_readdata                          => nios_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                               --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_nios_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_nios_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_nios_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_nios_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_nios_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_nios_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_nios_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_nios_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                -- custom_instruction_master.readra
		);

	pll : component PongFPGA_PLL
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_002_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_1_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_1_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_1_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_1_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_1_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => pll_c1_clk,                                --                    c1.clk
			c2                 => pll_c2_clk,                                --                    c2.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	vram : component PongFPGA_VRAM
		port map (
			clk         => pll_c0_clk,                             --   clk1.clk
			address     => mm_interconnect_1_vram_s1_address,      --     s1.address
			clken       => mm_interconnect_1_vram_s1_clken,        --       .clken
			chipselect  => mm_interconnect_1_vram_s1_chipselect,   --       .chipselect
			write       => mm_interconnect_1_vram_s1_write,        --       .write
			readdata    => mm_interconnect_1_vram_s1_readdata,     --       .readdata
			writedata   => mm_interconnect_1_vram_s1_writedata,    --       .writedata
			reset       => rst_controller_001_reset_out_reset,     -- reset1.reset
			reset_req   => rst_controller_001_reset_out_reset_req, --       .reset_req
			address2    => mm_interconnect_0_vram_s2_address,      --     s2.address
			chipselect2 => mm_interconnect_0_vram_s2_chipselect,   --       .chipselect
			clken2      => mm_interconnect_0_vram_s2_clken,        --       .clken
			write2      => mm_interconnect_0_vram_s2_write,        --       .write
			readdata2   => mm_interconnect_0_vram_s2_readdata,     --       .readdata
			writedata2  => mm_interconnect_0_vram_s2_writedata,    --       .writedata
			clk2        => pll_c1_clk,                             --   clk2.clk
			reset2      => rst_controller_reset_out_reset,         -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,     --       .reset_req
			freeze      => '0'                                     -- (terminated)
		);

	mm_interconnect_0 : component PongFPGA_mm_interconnect_0
		port map (
			PLL_c1_clk                                                     => pll_c1_clk,                                           --                                                   PLL_c1.clk
			AvalonRAMConnector_mono_1b_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- AvalonRAMConnector_mono_1b_0_reset_reset_bridge_in_reset.reset
			AvalonRAMConnector_mono_1b_0_avalon_master_address             => avalonramconnector_mono_1b_0_avalon_master_address,   --               AvalonRAMConnector_mono_1b_0_avalon_master.address
			AvalonRAMConnector_mono_1b_0_avalon_master_read                => avalonramconnector_mono_1b_0_avalon_master_read,      --                                                         .read
			AvalonRAMConnector_mono_1b_0_avalon_master_readdata            => avalonramconnector_mono_1b_0_avalon_master_readdata,  --                                                         .readdata
			AvalonRAMConnector_mono_1b_0_avalon_master_write               => avalonramconnector_mono_1b_0_avalon_master_write,     --                                                         .write
			AvalonRAMConnector_mono_1b_0_avalon_master_writedata           => avalonramconnector_mono_1b_0_avalon_master_writedata, --                                                         .writedata
			VRAM_s2_address                                                => mm_interconnect_0_vram_s2_address,                    --                                                  VRAM_s2.address
			VRAM_s2_write                                                  => mm_interconnect_0_vram_s2_write,                      --                                                         .write
			VRAM_s2_readdata                                               => mm_interconnect_0_vram_s2_readdata,                   --                                                         .readdata
			VRAM_s2_writedata                                              => mm_interconnect_0_vram_s2_writedata,                  --                                                         .writedata
			VRAM_s2_chipselect                                             => mm_interconnect_0_vram_s2_chipselect,                 --                                                         .chipselect
			VRAM_s2_clken                                                  => mm_interconnect_0_vram_s2_clken                       --                                                         .clken
		);

	mm_interconnect_1 : component PongFPGA_mm_interconnect_1
		port map (
			CLK_clk_clk                                           => clk_clk,                                            --                                         CLK_clk.clk
			PLL_c0_clk                                            => pll_c0_clk,                                         --                                          PLL_c0.clk
			NIOS_reset_reset_bridge_in_reset_reset                => rst_controller_001_reset_out_reset,                 --                NIOS_reset_reset_bridge_in_reset.reset
			PLL_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                 -- PLL_inclk_interface_reset_reset_bridge_in_reset.reset
			NIOS_data_master_address                              => nios_data_master_address,                           --                                NIOS_data_master.address
			NIOS_data_master_waitrequest                          => nios_data_master_waitrequest,                       --                                                .waitrequest
			NIOS_data_master_byteenable                           => nios_data_master_byteenable,                        --                                                .byteenable
			NIOS_data_master_read                                 => nios_data_master_read,                              --                                                .read
			NIOS_data_master_readdata                             => nios_data_master_readdata,                          --                                                .readdata
			NIOS_data_master_write                                => nios_data_master_write,                             --                                                .write
			NIOS_data_master_writedata                            => nios_data_master_writedata,                         --                                                .writedata
			NIOS_data_master_debugaccess                          => nios_data_master_debugaccess,                       --                                                .debugaccess
			NIOS_instruction_master_address                       => nios_instruction_master_address,                    --                         NIOS_instruction_master.address
			NIOS_instruction_master_waitrequest                   => nios_instruction_master_waitrequest,                --                                                .waitrequest
			NIOS_instruction_master_read                          => nios_instruction_master_read,                       --                                                .read
			NIOS_instruction_master_readdata                      => nios_instruction_master_readdata,                   --                                                .readdata
			NIOS_debug_mem_slave_address                          => mm_interconnect_1_nios_debug_mem_slave_address,     --                            NIOS_debug_mem_slave.address
			NIOS_debug_mem_slave_write                            => mm_interconnect_1_nios_debug_mem_slave_write,       --                                                .write
			NIOS_debug_mem_slave_read                             => mm_interconnect_1_nios_debug_mem_slave_read,        --                                                .read
			NIOS_debug_mem_slave_readdata                         => mm_interconnect_1_nios_debug_mem_slave_readdata,    --                                                .readdata
			NIOS_debug_mem_slave_writedata                        => mm_interconnect_1_nios_debug_mem_slave_writedata,   --                                                .writedata
			NIOS_debug_mem_slave_byteenable                       => mm_interconnect_1_nios_debug_mem_slave_byteenable,  --                                                .byteenable
			NIOS_debug_mem_slave_waitrequest                      => mm_interconnect_1_nios_debug_mem_slave_waitrequest, --                                                .waitrequest
			NIOS_debug_mem_slave_debugaccess                      => mm_interconnect_1_nios_debug_mem_slave_debugaccess, --                                                .debugaccess
			PLL_pll_slave_address                                 => mm_interconnect_1_pll_pll_slave_address,            --                                   PLL_pll_slave.address
			PLL_pll_slave_write                                   => mm_interconnect_1_pll_pll_slave_write,              --                                                .write
			PLL_pll_slave_read                                    => mm_interconnect_1_pll_pll_slave_read,               --                                                .read
			PLL_pll_slave_readdata                                => mm_interconnect_1_pll_pll_slave_readdata,           --                                                .readdata
			PLL_pll_slave_writedata                               => mm_interconnect_1_pll_pll_slave_writedata,          --                                                .writedata
			VRAM_s1_address                                       => mm_interconnect_1_vram_s1_address,                  --                                         VRAM_s1.address
			VRAM_s1_write                                         => mm_interconnect_1_vram_s1_write,                    --                                                .write
			VRAM_s1_readdata                                      => mm_interconnect_1_vram_s1_readdata,                 --                                                .readdata
			VRAM_s1_writedata                                     => mm_interconnect_1_vram_s1_writedata,                --                                                .writedata
			VRAM_s1_chipselect                                    => mm_interconnect_1_vram_s1_chipselect,               --                                                .chipselect
			VRAM_s1_clken                                         => mm_interconnect_1_vram_s1_clken                     --                                                .clken
		);

	irq_mapper : component PongFPGA_irq_mapper
		port map (
			clk        => pll_c0_clk,                         --       clk.clk
			reset      => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sender_irq => nios_irq_irq                        --    sender.irq
		);

	rst_controller : component pongfpga_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_c1_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component pongfpga_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => pll_c0_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component pongfpga_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of PongFPGA
