-- PongFPGA.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PongFPGA is
	port (
		clk_clk                     : in  std_logic                    := '0'; --             clk.clk
		hdmidriver_hdmi_output_clk  : out std_logic;                           -- hdmidriver_hdmi.output_clk
		hdmidriver_hdmi_output_data : out std_logic_vector(2 downto 0);        --                .output_data
		reset_reset_n               : in  std_logic                    := '0'  --           reset.reset_n
	);
end entity PongFPGA;

architecture rtl of PongFPGA is
	component HDMIDriver is
		generic (
			DISPLAY_RES_WIDTH  : integer := 640;
			DISPLAY_RES_HEIGHT : integer := 480;
			PX_FRONT_PORCH     : integer := 16;
			PX_SYNC_PULSE      : integer := 96;
			PX_BACK_PORCH      : integer := 48;
			ROW_FRONT_PORCH    : integer := 10;
			ROW_SYNC_PULSE     : integer := 2;
			ROW_BACK_PORCH     : integer := 33
		);
		port (
			clk         : in  std_logic                     := 'X'; -- clk
			HDMI_clk    : in  std_logic                     := 'X'; -- clk
			output_clk  : out std_logic;                            -- output_clk
			output_data : out std_logic_vector(2 downto 0);         -- output_data
			px_color    : in  std_logic                     := 'X'; -- px_color
			px_x        : out std_logic_vector(12 downto 0);        -- px_x
			px_y        : out std_logic_vector(12 downto 0)         -- px_y
		);
	end component HDMIDriver;

	component HDMIImageGenerator is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			px_color : out std_logic;                                        -- px_color
			px_x     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- px_x
			px_y     : in  std_logic_vector(12 downto 0) := (others => 'X')  -- px_y
		);
	end component HDMIImageGenerator;

	component PongFPGA_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component PongFPGA_altpll_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal altpll_0_c0_clk                                      : std_logic;                     -- altpll_0:c0 -> [HDMIDriver_0:clk, HDMI_IMAGE_GEN_MONO_1b_0:clk]
	signal altpll_0_c1_clk                                      : std_logic;                     -- altpll_0:c1 -> HDMIDriver_0:HDMI_clk
	signal hdmidriver_0_px_address_px_x                         : std_logic_vector(12 downto 0); -- HDMIDriver_0:px_x -> HDMI_IMAGE_GEN_MONO_1b_0:px_x
	signal hdmidriver_0_px_address_px_y                         : std_logic_vector(12 downto 0); -- HDMIDriver_0:px_y -> HDMI_IMAGE_GEN_MONO_1b_0:px_y
	signal hdmi_image_gen_mono_1b_0_hdmiimagegenerator_px_color : std_logic;                     -- HDMI_IMAGE_GEN_MONO_1b_0:px_color -> HDMIDriver_0:px_color
	signal altpll_0_locked_conduit_export                       : std_logic;                     -- altpll_0:locked -> altpll_0:areset
	signal rst_controller_reset_out_reset                       : std_logic;                     -- rst_controller:reset_out -> altpll_0:reset
	signal reset_reset_n_ports_inv                              : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	hdmidriver_0 : component HDMIDriver
		generic map (
			DISPLAY_RES_WIDTH  => 640,
			DISPLAY_RES_HEIGHT => 480,
			PX_FRONT_PORCH     => 16,
			PX_SYNC_PULSE      => 96,
			PX_BACK_PORCH      => 48,
			ROW_FRONT_PORCH    => 10,
			ROW_SYNC_PULSE     => 2,
			ROW_BACK_PORCH     => 33
		)
		port map (
			clk         => altpll_0_c0_clk,                                      --      clock.clk
			HDMI_clk    => altpll_0_c1_clk,                                      --   HDMI_clk.clk
			output_clk  => hdmidriver_hdmi_output_clk,                           --       HDMI.output_clk
			output_data => hdmidriver_hdmi_output_data,                          --           .output_data
			px_color    => hdmi_image_gen_mono_1b_0_hdmiimagegenerator_px_color, --   PX_COLOR.px_color
			px_x        => hdmidriver_0_px_address_px_x,                         -- PX_ADDRESS.px_x
			px_y        => hdmidriver_0_px_address_px_y                          --           .px_y
		);

	hdmi_image_gen_mono_1b_0 : component HDMIImageGenerator
		port map (
			clk      => altpll_0_c0_clk,                                      --              clock.clk
			px_color => hdmi_image_gen_mono_1b_0_hdmiimagegenerator_px_color, -- HDMIImageGenerator.px_color
			px_x     => hdmidriver_0_px_address_px_x,                         --         PX_ADDRESS.px_x
			px_y     => hdmidriver_0_px_address_px_y                          --                   .px_y
		);

	altpll_0 : component PongFPGA_altpll_0
		port map (
			clk                => clk_clk,                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset, -- inclk_interface_reset.reset
			read               => open,                           --             pll_slave.read
			write              => open,                           --                      .write
			address            => open,                           --                      .address
			readdata           => open,                           --                      .readdata
			writedata          => open,                           --                      .writedata
			c0                 => altpll_0_c0_clk,                --                    c0.clk
			c1                 => altpll_0_c1_clk,                --                    c1.clk
			areset             => altpll_0_locked_conduit_export, --        areset_conduit.export
			locked             => altpll_0_locked_conduit_export, --        locked_conduit.export
			scandone           => open,                           --           (terminated)
			scandataout        => open,                           --           (terminated)
			c2                 => open,                           --           (terminated)
			c3                 => open,                           --           (terminated)
			c4                 => open,                           --           (terminated)
			phasedone          => open,                           --           (terminated)
			phasecounterselect => "000",                          --           (terminated)
			phaseupdown        => '0',                            --           (terminated)
			phasestep          => '0',                            --           (terminated)
			scanclk            => '0',                            --           (terminated)
			scanclkena         => '0',                            --           (terminated)
			scandata           => '0',                            --           (terminated)
			configupdate       => '0'                             --           (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of PongFPGA
