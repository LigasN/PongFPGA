-- PongFPGA_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PongFPGA_tb is
end entity PongFPGA_tb;

architecture rtl of PongFPGA_tb is
	component PongFPGA is
		port (
			clk_clk                     : in  std_logic                    := 'X'; -- clk
			hdmidriver_hdmi_output_clk  : out std_logic;                           -- output_clk
			hdmidriver_hdmi_output_data : out std_logic_vector(2 downto 0);        -- output_data
			reset_reset_n               : in  std_logic                    := 'X'  -- reset_n
		);
	end component PongFPGA;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			clk             : in std_logic                    := 'X';             -- clk
			sig_output_clk  : in std_logic_vector(0 downto 0) := (others => 'X'); -- output_clk
			sig_output_data : in std_logic_vector(2 downto 0) := (others => 'X'); -- output_data
			reset           : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal pongfpga_inst_clk_bfm_clk_clk             : std_logic;                    -- PongFPGA_inst_clk_bfm:clk -> [PongFPGA_inst:clk_clk, PongFPGA_inst_hdmidriver_hdmi_bfm:clk, PongFPGA_inst_reset_bfm:clk]
	signal pongfpga_inst_hdmidriver_hdmi_output_clk  : std_logic;                    -- PongFPGA_inst:hdmidriver_hdmi_output_clk -> PongFPGA_inst_hdmidriver_hdmi_bfm:sig_output_clk
	signal pongfpga_inst_hdmidriver_hdmi_output_data : std_logic_vector(2 downto 0); -- PongFPGA_inst:hdmidriver_hdmi_output_data -> PongFPGA_inst_hdmidriver_hdmi_bfm:sig_output_data
	signal pongfpga_inst_reset_bfm_reset_reset       : std_logic;                    -- PongFPGA_inst_reset_bfm:reset -> PongFPGA_inst:reset_reset_n

begin

	pongfpga_inst : component PongFPGA
		port map (
			clk_clk                     => pongfpga_inst_clk_bfm_clk_clk,             --             clk.clk
			hdmidriver_hdmi_output_clk  => pongfpga_inst_hdmidriver_hdmi_output_clk,  -- hdmidriver_hdmi.output_clk
			hdmidriver_hdmi_output_data => pongfpga_inst_hdmidriver_hdmi_output_data, --                .output_data
			reset_reset_n               => pongfpga_inst_reset_bfm_reset_reset        --           reset.reset_n
		);

	pongfpga_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 10000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => pongfpga_inst_clk_bfm_clk_clk  -- clk.clk
		);

	pongfpga_inst_hdmidriver_hdmi_bfm : component altera_conduit_bfm
		port map (
			clk               => pongfpga_inst_clk_bfm_clk_clk,             --     clk.clk
			sig_output_clk(0) => pongfpga_inst_hdmidriver_hdmi_output_clk,  -- conduit.output_clk
			sig_output_data   => pongfpga_inst_hdmidriver_hdmi_output_data, --        .output_data
			reset             => '0'                                        -- (terminated)
		);

	pongfpga_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => pongfpga_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => pongfpga_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of PongFPGA_tb
